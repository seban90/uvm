`define AXI_FIXED 2'b00
`define AXI_INCR  2'b01
`define AXI_WRAP  2'b10

`define AXI_1_BYTE   3'b000
`define AXI_2_BYTE   3'b001
`define AXI_4_BYTE   3'b010
`define AXI_8_BYTE   3'b011
`define AXI_16_BYTE  3'b100
`define AXI_32_BYTE  3'b101
`define AXI_64_BYTE  3'b110
`define AXI_128_BYTE 3'b111
